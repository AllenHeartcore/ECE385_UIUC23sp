module FontROM (
	input  logic [10:0] addr,
	output logic [ 7:0] data);

	parameter ADDR_WIDTH = 11;
	parameter DATA_WIDTH =  8;

	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7E, 8'h81, 8'hA5, 8'h81, 8'h81, 8'hBD, 8'h99, 8'h81, 8'h81, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7E, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hC3, 8'hE7, 8'hFF, 8'hFF, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h6C, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'h7C, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h38, 8'h7C, 8'hFE, 8'h7C, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'hE7, 8'hE7, 8'hE7, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'hFF, 8'hFF, 8'h7E, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hC3, 8'hC3, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h66, 8'h42, 8'h42, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h99, 8'hBD, 8'hBD, 8'h99, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
	8'h00, 8'h00, 8'h1E, 8'h0E, 8'h1A, 8'h32, 8'h78, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h18, 8'h7E, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3F, 8'h33, 8'h3F, 8'h30, 8'h30, 8'h30, 8'h30, 8'h70, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7F, 8'h63, 8'h7F, 8'h63, 8'h63, 8'h63, 8'h63, 8'h67, 8'hE7, 8'hE6, 8'hC0, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'hDB, 8'h3C, 8'hE7, 8'h3C, 8'hDB, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h80, 8'hC0, 8'hE0, 8'hF0, 8'hF8, 8'hFE, 8'hF8, 8'hF0, 8'hE0, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h02, 8'h06, 8'h0E, 8'h1E, 8'h3E, 8'hFE, 8'h3E, 8'h1E, 8'h0E, 8'h06, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h00, 8'h66, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7F, 8'hDB, 8'hDB, 8'hDB, 8'h7B, 8'h1B, 8'h1B, 8'h1B, 8'h1B, 8'h1B, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h7C, 8'hC6, 8'h60, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'h6C, 8'h38, 8'h0C, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h0C, 8'hFE, 8'h0C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h60, 8'hFE, 8'h60, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hC0, 8'hC0, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h66, 8'hFF, 8'h66, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h38, 8'h38, 8'h7C, 8'h7C, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'h7C, 8'h7C, 8'h38, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h66, 8'h66, 8'h66, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h6C, 8'h6C, 8'hFE, 8'h6C, 8'h6C, 8'h6C, 8'hFE, 8'h6C, 8'h6C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h18, 8'h18, 8'h7C, 8'hC6, 8'hC2, 8'hC0, 8'h7C, 8'h06, 8'h06, 8'h86, 8'hC6, 8'h7C, 8'h18, 8'h18, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'hC2, 8'hC6, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC6, 8'h86, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h6C, 8'h6C, 8'h38, 8'h76, 8'hDC, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h30, 8'h30, 8'h30, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h0C, 8'h18, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h18, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h30, 8'h18, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h66, 8'h3C, 8'hFF, 8'h3C, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h7E, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hCE, 8'hDE, 8'hF6, 8'hE6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h38, 8'h78, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC0, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'h06, 8'h06, 8'h3C, 8'h06, 8'h06, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h0C, 8'h1C, 8'h3C, 8'h6C, 8'hCC, 8'hFE, 8'h0C, 8'h0C, 8'h0C, 8'h1E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'hC0, 8'hC0, 8'hC0, 8'hFC, 8'h06, 8'h06, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h60, 8'hC0, 8'hC0, 8'hFC, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'hC6, 8'h06, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h30, 8'h30, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'h7E, 8'h06, 8'h06, 8'h06, 8'h0C, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'h0C, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hDE, 8'hDE, 8'hDE, 8'hDC, 8'hC0, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h10, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFC, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h66, 8'h66, 8'h66, 8'h66, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h66, 8'hC2, 8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hC2, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hF8, 8'h6C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h6C, 8'hF8, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'h66, 8'h62, 8'h68, 8'h78, 8'h68, 8'h60, 8'h62, 8'h66, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'h66, 8'h62, 8'h68, 8'h78, 8'h68, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h66, 8'hC2, 8'hC0, 8'hC0, 8'hDE, 8'hC6, 8'hC6, 8'h66, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h1E, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'hCC, 8'hCC, 8'hCC, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hE6, 8'h66, 8'h66, 8'h6C, 8'h78, 8'h78, 8'h6C, 8'h66, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hF0, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h62, 8'h66, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hE7, 8'hFF, 8'hFF, 8'hDB, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC6, 8'hE6, 8'hF6, 8'hFE, 8'hDE, 8'hCE, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFC, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h60, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hD6, 8'hDE, 8'h7C, 8'h0C, 8'h0E, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFC, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h6C, 8'h66, 8'h66, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'h60, 8'h38, 8'h0C, 8'h06, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFF, 8'hDB, 8'h99, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hDB, 8'hDB, 8'hFF, 8'h66, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h3C, 8'h66, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFF, 8'hC3, 8'h86, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC1, 8'hC3, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h80, 8'hC0, 8'hE0, 8'h70, 8'h38, 8'h1C, 8'h0E, 8'h06, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h10, 8'h38, 8'h6C, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00,
	8'h30, 8'h30, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h78, 8'h0C, 8'h7C, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hE0, 8'h60, 8'h60, 8'h78, 8'h6C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC0, 8'hC0, 8'hC0, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h1C, 8'h0C, 8'h0C, 8'h3C, 8'h6C, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'hFE, 8'hC0, 8'hC0, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h6C, 8'h64, 8'h60, 8'hF0, 8'h60, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h76, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h7C, 8'h0C, 8'hCC, 8'h78, 8'h00,
	8'h00, 8'h00, 8'hE0, 8'h60, 8'h60, 8'h6C, 8'h76, 8'h66, 8'h66, 8'h66, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h06, 8'h06, 8'h00, 8'h0E, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h66, 8'h66, 8'h3C, 8'h00,
	8'h00, 8'h00, 8'hE0, 8'h60, 8'h60, 8'h66, 8'h6C, 8'h78, 8'h78, 8'h6C, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hE6, 8'hFF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDC, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDC, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h60, 8'h60, 8'hF0, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h76, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h7C, 8'h0C, 8'h0C, 8'h1E, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDC, 8'h76, 8'h66, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'h60, 8'h38, 8'h0C, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h10, 8'h30, 8'h30, 8'hFC, 8'h30, 8'h30, 8'h30, 8'h30, 8'h36, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hDB, 8'hDB, 8'hFF, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h3C, 8'h66, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7E, 8'h06, 8'h0C, 8'hF8, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hCC, 8'h18, 8'h30, 8'h60, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h0E, 8'h18, 8'h18, 8'h18, 8'h70, 8'h18, 8'h18, 8'h18, 8'h18, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h70, 8'h18, 8'h18, 8'h18, 8'h0E, 8'h18, 8'h18, 8'h18, 8'h18, 8'h70, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};

	assign data = ROM[addr];

endmodule
