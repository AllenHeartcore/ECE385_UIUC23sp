module I2S (
	input  logic SCLK, LRCLK, DIN,
	output logic DOUT);


endmodule
