/* [MapROM Entry Format]
 * |     19-14      |      13-6      |  5-0   |
 * | DrawYAnch[9:4] | DrawXAnch[9:2] | keyidx |
 *
 * Each entry encodes the region assignment of a 56x4 block.
 *
 * [keyidx (keycode - 5) Positions]
 * 26  27  28  29  30  31  32  33  34  40  41
 *   21   3  16  18  23  19   7  13  14  42
 *     17   2   4   5   6   8   9  10  46
 *       22   1  20   0  12  11  49  50
 */


module MapROM (
	input  logic [ 9:0] addr,
	output logic [19:0] data);

	parameter [0:639][19:0] ROM = {
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA,
	20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA, 20'h400DA,
	20'h400DA, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B,
	20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h4045B, 20'h407DC,
	20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC,
	20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC, 20'h407DC, 20'h40B5D, 20'h40B5D, 20'h40B5D,
	20'h40B5D, 20'h40B5D, 20'h40B5D, 20'h40B5D, 20'h40B5D, 20'h40B5D, 20'h40B5D, 20'h40B5D,
	20'h40B5D, 20'h40B5D, 20'h40B5D, 20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE,
	20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE, 20'h40EDE,
	20'h40EDE, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F,
	20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h4125F, 20'h415E0,
	20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0,
	20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0, 20'h415E0, 20'h41961, 20'h41961, 20'h41961,
	20'h41961, 20'h41961, 20'h41961, 20'h41961, 20'h41961, 20'h41961, 20'h41961, 20'h41961,
	20'h41961, 20'h41961, 20'h41961, 20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2,
	20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2, 20'h41CE2,
	20'h41CE2, 20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h42068,
	20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h42068, 20'h423E9,
	20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9,
	20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9, 20'h423E9, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295,
	20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295, 20'h5C295,
	20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603,
	20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C603, 20'h5C990, 20'h5C990,
	20'h5C990, 20'h5C990, 20'h5C990, 20'h5C990, 20'h5C990, 20'h5C990, 20'h5C990, 20'h5C990,
	20'h5C990, 20'h5C990, 20'h5C990, 20'h5C990, 20'h5CD12, 20'h5CD12, 20'h5CD12, 20'h5CD12,
	20'h5CD12, 20'h5CD12, 20'h5CD12, 20'h5CD12, 20'h5CD12, 20'h5CD12, 20'h5CD12, 20'h5CD12,
	20'h5CD12, 20'h5CD12, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097,
	20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097, 20'h5D097,
	20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413,
	20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D413, 20'h5D787, 20'h5D787,
	20'h5D787, 20'h5D787, 20'h5D787, 20'h5D787, 20'h5D787, 20'h5D787, 20'h5D787, 20'h5D787,
	20'h5D787, 20'h5D787, 20'h5D787, 20'h5D787, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D,
	20'h5DB0D, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D, 20'h5DB0D,
	20'h5DB0D, 20'h5DB0D, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E,
	20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E, 20'h5DE8E,
	20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A,
	20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'h5E22A, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h78451,
	20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h78451, 20'h787C2,
	20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2,
	20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2, 20'h787C2, 20'h78B44, 20'h78B44, 20'h78B44,
	20'h78B44, 20'h78B44, 20'h78B44, 20'h78B44, 20'h78B44, 20'h78B44, 20'h78B44, 20'h78B44,
	20'h78B44, 20'h78B44, 20'h78B44, 20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5,
	20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5, 20'h78EC5,
	20'h78EC5, 20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h79246,
	20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h79246, 20'h795C8,
	20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8,
	20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8, 20'h795C8, 20'h79949, 20'h79949, 20'h79949,
	20'h79949, 20'h79949, 20'h79949, 20'h79949, 20'h79949, 20'h79949, 20'h79949, 20'h79949,
	20'h79949, 20'h79949, 20'h79949, 20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA,
	20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA, 20'h79CCA,
	20'h79CCA, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E,
	20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'h7A06E, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94616,
	20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94616, 20'h94981, 20'h94981,
	20'h94981, 20'h94981, 20'h94981, 20'h94981, 20'h94981, 20'h94981, 20'h94981, 20'h94981,
	20'h94981, 20'h94981, 20'h94981, 20'h94981, 20'h94D14, 20'h94D14, 20'h94D14, 20'h94D14,
	20'h94D14, 20'h94D14, 20'h94D14, 20'h94D14, 20'h94D14, 20'h94D14, 20'h94D14, 20'h94D14,
	20'h94D14, 20'h94D14, 20'h95080, 20'h95080, 20'h95080, 20'h95080, 20'h95080, 20'h95080,
	20'h95080, 20'h95080, 20'h95080, 20'h95080, 20'h95080, 20'h95080, 20'h95080, 20'h95080,
	20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C,
	20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9540C, 20'h9578B, 20'h9578B,
	20'h9578B, 20'h9578B, 20'h9578B, 20'h9578B, 20'h9578B, 20'h9578B, 20'h9578B, 20'h9578B,
	20'h9578B, 20'h9578B, 20'h9578B, 20'h9578B, 20'h95B31, 20'h95B31, 20'h95B31, 20'h95B31,
	20'h95B31, 20'h95B31, 20'h95B31, 20'h95B31, 20'h95B31, 20'h95B31, 20'h95B31, 20'h95B31,
	20'h95B31, 20'h95B31, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2,
	20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2, 20'h95EB2,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF,
	20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF, 20'hFFFFF};

	assign data = ROM[addr];

endmodule


module FontROM (
	input  logic [10:0] addr,
	output logic [ 7:0] data);

	parameter ADDR_WIDTH = 11;
	parameter DATA_WIDTH =  8;

	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7E, 8'h81, 8'hA5, 8'h81, 8'h81, 8'hBD, 8'h99, 8'h81, 8'h81, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7E, 8'hFF, 8'hDB, 8'hFF, 8'hFF, 8'hC3, 8'hE7, 8'hFF, 8'hFF, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h6C, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'h7C, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h38, 8'h7C, 8'hFE, 8'h7C, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'hE7, 8'hE7, 8'hE7, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'hFF, 8'hFF, 8'h7E, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hC3, 8'hC3, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h66, 8'h42, 8'h42, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h99, 8'hBD, 8'hBD, 8'h99, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
	8'h00, 8'h00, 8'h1E, 8'h0E, 8'h1A, 8'h32, 8'h78, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h3C, 8'h18, 8'h7E, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3F, 8'h33, 8'h3F, 8'h30, 8'h30, 8'h30, 8'h30, 8'h70, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7F, 8'h63, 8'h7F, 8'h63, 8'h63, 8'h63, 8'h63, 8'h67, 8'hE7, 8'hE6, 8'hC0, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'hDB, 8'h3C, 8'hE7, 8'h3C, 8'hDB, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h80, 8'hC0, 8'hE0, 8'hF0, 8'hF8, 8'hFE, 8'hF8, 8'hF0, 8'hE0, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h02, 8'h06, 8'h0E, 8'h1E, 8'h3E, 8'hFE, 8'h3E, 8'h1E, 8'h0E, 8'h06, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h00, 8'h66, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7F, 8'hDB, 8'hDB, 8'hDB, 8'h7B, 8'h1B, 8'h1B, 8'h1B, 8'h1B, 8'h1B, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h7C, 8'hC6, 8'h60, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'h6C, 8'h38, 8'h0C, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h7E, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h0C, 8'hFE, 8'h0C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h60, 8'hFE, 8'h60, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hC0, 8'hC0, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h66, 8'hFF, 8'h66, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h38, 8'h38, 8'h7C, 8'h7C, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'h7C, 8'h7C, 8'h38, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h66, 8'h66, 8'h66, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h6C, 8'h6C, 8'hFE, 8'h6C, 8'h6C, 8'h6C, 8'hFE, 8'h6C, 8'h6C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h18, 8'h18, 8'h7C, 8'hC6, 8'hC2, 8'hC0, 8'h7C, 8'h06, 8'h06, 8'h86, 8'hC6, 8'h7C, 8'h18, 8'h18, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'hC2, 8'hC6, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC6, 8'h86, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h6C, 8'h6C, 8'h38, 8'h76, 8'hDC, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h30, 8'h30, 8'h30, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h0C, 8'h18, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h18, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h30, 8'h18, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h66, 8'h3C, 8'hFF, 8'h3C, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h7E, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hCE, 8'hDE, 8'hF6, 8'hE6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h38, 8'h78, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC0, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'h06, 8'h06, 8'h3C, 8'h06, 8'h06, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h0C, 8'h1C, 8'h3C, 8'h6C, 8'hCC, 8'hFE, 8'h0C, 8'h0C, 8'h0C, 8'h1E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'hC0, 8'hC0, 8'hC0, 8'hFC, 8'h06, 8'h06, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h60, 8'hC0, 8'hC0, 8'hFC, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'hC6, 8'h06, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h30, 8'h30, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'h7E, 8'h06, 8'h06, 8'h06, 8'h0C, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h60, 8'h30, 8'h18, 8'h0C, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'h0C, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hDE, 8'hDE, 8'hDE, 8'hDC, 8'hC0, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h10, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFC, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h66, 8'h66, 8'h66, 8'h66, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h66, 8'hC2, 8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hC2, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hF8, 8'h6C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h6C, 8'hF8, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'h66, 8'h62, 8'h68, 8'h78, 8'h68, 8'h60, 8'h62, 8'h66, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFE, 8'h66, 8'h62, 8'h68, 8'h78, 8'h68, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h66, 8'hC2, 8'hC0, 8'hC0, 8'hDE, 8'hC6, 8'hC6, 8'h66, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h1E, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'hCC, 8'hCC, 8'hCC, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hE6, 8'h66, 8'h66, 8'h6C, 8'h78, 8'h78, 8'h6C, 8'h66, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hF0, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h62, 8'h66, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hE7, 8'hFF, 8'hFF, 8'hDB, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC6, 8'hE6, 8'hF6, 8'hFE, 8'hDE, 8'hCE, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFC, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h60, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hD6, 8'hDE, 8'h7C, 8'h0C, 8'h0E, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFC, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h6C, 8'h66, 8'h66, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'h60, 8'h38, 8'h0C, 8'h06, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFF, 8'hDB, 8'h99, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'hDB, 8'hDB, 8'hFF, 8'h66, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h3C, 8'h66, 8'hC3, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hFF, 8'hC3, 8'h86, 8'h0C, 8'h18, 8'h30, 8'h60, 8'hC1, 8'hC3, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h30, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h80, 8'hC0, 8'hE0, 8'h70, 8'h38, 8'h1C, 8'h0E, 8'h06, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h3C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h10, 8'h38, 8'h6C, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00,
	8'h30, 8'h30, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h78, 8'h0C, 8'h7C, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'hE0, 8'h60, 8'h60, 8'h78, 8'h6C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC0, 8'hC0, 8'hC0, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h1C, 8'h0C, 8'h0C, 8'h3C, 8'h6C, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'hFE, 8'hC0, 8'hC0, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h6C, 8'h64, 8'h60, 8'hF0, 8'h60, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h76, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h7C, 8'h0C, 8'hCC, 8'h78, 8'h00,
	8'h00, 8'h00, 8'hE0, 8'h60, 8'h60, 8'h6C, 8'h76, 8'h66, 8'h66, 8'h66, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h18, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h06, 8'h06, 8'h00, 8'h0E, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h66, 8'h66, 8'h3C, 8'h00,
	8'h00, 8'h00, 8'hE0, 8'h60, 8'h60, 8'h66, 8'h6C, 8'h78, 8'h78, 8'h6C, 8'h66, 8'hE6, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hE6, 8'hFF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDC, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDC, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h7C, 8'h60, 8'h60, 8'hF0, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h76, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h7C, 8'h0C, 8'h0C, 8'h1E, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDC, 8'h76, 8'h66, 8'h60, 8'h60, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hC6, 8'h60, 8'h38, 8'h0C, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h10, 8'h30, 8'h30, 8'hFC, 8'h30, 8'h30, 8'h30, 8'h30, 8'h36, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h76, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'hC3, 8'hC3, 8'hDB, 8'hDB, 8'hFF, 8'h66, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'h66, 8'h3C, 8'h18, 8'h3C, 8'h66, 8'hC3, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7E, 8'h06, 8'h0C, 8'hF8, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hCC, 8'h18, 8'h30, 8'h60, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h0E, 8'h18, 8'h18, 8'h18, 8'h70, 8'h18, 8'h18, 8'h18, 8'h18, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h70, 8'h18, 8'h18, 8'h18, 8'h0E, 8'h18, 8'h18, 8'h18, 8'h18, 8'h70, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h76, 8'hDC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
	8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hC6, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};

	assign data = ROM[addr];

endmodule
